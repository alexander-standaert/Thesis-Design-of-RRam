.SUBCKT memristor_ieee Pos Neg PARAM:

*Parameters:
n=4 a1=9 a2=0.01 b1=2 b2=4 l=10n
wmin=0.05 wmax=0.95 p0=1.2 fon=40E-3 foff=40E-3

*Shape facor, sf, can be a function of tunneling barrier width (normalized state variable)
sfo=4 sfm=20 p=5 *** sf(w)=sfo+sfm(1-(2w)**2p)

*State variable:
Gvon 0 w value = signm(wmax-V(w))*signm(V(Pos,Neg))*gon(V(Pos,Neg),sf(V(w)),po)
Gvoff 0 w value = signm(V(w)-wmin)*signm(V(Neg,Pos))*goff(V(Pos,Neg),sf(V(w)),p0)

*Initial (internal) state:
.IC V(w) 0.5

*Integration:
Cw w 0 8e-5
Rw w 0 0.01T

*Current equation:
Gmem Pos Neg value = l*((V(w)**n)*a1*sinh(b1*V(Pos,Neg))+a2*(exp(b2*V(Pos,Neg))-1))

*Series resistor Rs, can be implemented here, between two Neg1 and Neg2 nodes.

*Functions:
.func signm(v) = (sgn(v)+1)/2
.func gon(v1,v2,v3) = fon*((1-v1/(2*v3))*exp(v2*v3*(1-sqrt((1-v1/(2*v3))))))
.func goff(v1,v2,v3) = foff*(-((1+v1/(2*v3))*exp(v2*v3*(1-sqrt((1+v1/(2*v3)))))))
.func sf(v1) = sfo+sfm(1-(2*(v1)-1)**2p)

.END memristor_ieee
