* hspice / eldo example

* --------------------------------
* needed for eldo :
.PROBE DC
.PROBE TRAN
* ------------------------------

.OPTIONS CSDF

.TRAN 0.1p  10n
.DC Vin 0 1 0.1

* to generate the netlist: use:
* mat2spice( 'RClong.m2s', 'generatedNetlist' )

Vin n1 0 pulse 0 1 1n 0.1n 0.2n 0.4n 1n 
*Vin  n1 0 PWL( 0p 0 10p 1 )

R_1   n2 n1 1
C_1   n2 0      1f

R_2   n3 n2 1
C_2   n3 0      1f

R_3   n4 n3 1
C_3   n4 0      1f

R_4   n5 n4 1
C_4   n5 0      1f

R_5   n6 n5 1
C_5   n6 0      1f

R_6   n7 n6 1
C_6   n7 0      1f

R_7   n8 n7 1
C_7   n8 0      1f

R_8   n9 n8 1
C_8   n9 0      1f

R_9   n10 n9 1
C_9   n10 0      1f

R_10   n11 n10 1
C_10   n11 0      1f

R_11   n12 n11 1
C_11   n12 0      1f

R_12   n13 n12 1
C_12   n13 0      1f

R_13   n14 n13 1
C_13   n14 0      1f

R_14   n15 n14 1
C_14   n15 0      1f

R_15   n16 n15 1
C_15   n16 0      1f

R_16   n17 n16 1
C_16   n17 0      1f

R_17   n18 n17 1
C_17   n18 0      1f

R_18   n19 n18 1
C_18   n19 0      1f

R_19   n20 n19 1
C_19   n20 0      1f

R_20   n21 n20 1
C_20   n21 0      1f

R_21   n22 n21 1
C_21   n22 0      1f

R_22   n23 n22 1
C_22   n23 0      1f

R_23   n24 n23 1
C_23   n24 0      1f

R_24   n25 n24 1
C_24   n25 0      1f

R_25   n26 n25 1
C_25   n26 0      1f

R_26   n27 n26 1
C_26   n27 0      1f

R_27   n28 n27 1
C_27   n28 0      1f

R_28   n29 n28 1
C_28   n29 0      1f

R_29   n30 n29 1
C_29   n30 0      1f

R_30   n31 n30 1
C_30   n31 0      1f

R_31   n32 n31 1
C_31   n32 0      1f

R_32   n33 n32 1
C_32   n33 0      1f

R_33   n34 n33 1
C_33   n34 0      1f

R_34   n35 n34 1
C_34   n35 0      1f

R_35   n36 n35 1
C_35   n36 0      1f

R_36   n37 n36 1
C_36   n37 0      1f

R_37   n38 n37 1
C_37   n38 0      1f

R_38   n39 n38 1
C_38   n39 0      1f

R_39   n40 n39 1
C_39   n40 0      1f

R_40   n41 n40 1
C_40   n41 0      1f

R_41   n42 n41 1
C_41   n42 0      1f

R_42   n43 n42 1
C_42   n43 0      1f

R_43   n44 n43 1
C_43   n44 0      1f

R_44   n45 n44 1
C_44   n45 0      1f

R_45   n46 n45 1
C_45   n46 0      1f

R_46   n47 n46 1
C_46   n47 0      1f

R_47   n48 n47 1
C_47   n48 0      1f

R_48   n49 n48 1
C_48   n49 0      1f

R_49   n50 n49 1
C_49   n50 0      1f

R_50   n51 n50 1
C_50   n51 0      1f

R_51   n52 n51 1
C_51   n52 0      1f

R_52   n53 n52 1
C_52   n53 0      1f

R_53   n54 n53 1
C_53   n54 0      1f

R_54   n55 n54 1
C_54   n55 0      1f

R_55   n56 n55 1
C_55   n56 0      1f

R_56   n57 n56 1
C_56   n57 0      1f

R_57   n58 n57 1
C_57   n58 0      1f

R_58   n59 n58 1
C_58   n59 0      1f

R_59   n60 n59 1
C_59   n60 0      1f

R_60   n61 n60 1
C_60   n61 0      1f

R_61   n62 n61 1
C_61   n62 0      1f

R_62   n63 n62 1
C_62   n63 0      1f

R_63   n64 n63 1
C_63   n64 0      1f

R_64   n65 n64 1
C_64   n65 0      1f

R_65   n66 n65 1
C_65   n66 0      1f

R_66   n67 n66 1
C_66   n67 0      1f

R_67   n68 n67 1
C_67   n68 0      1f

R_68   n69 n68 1
C_68   n69 0      1f

R_69   n70 n69 1
C_69   n70 0      1f

R_70   n71 n70 1
C_70   n71 0      1f

R_71   n72 n71 1
C_71   n72 0      1f

R_72   n73 n72 1
C_72   n73 0      1f

R_73   n74 n73 1
C_73   n74 0      1f

R_74   n75 n74 1
C_74   n75 0      1f

R_75   n76 n75 1
C_75   n76 0      1f

R_76   n77 n76 1
C_76   n77 0      1f

R_77   n78 n77 1
C_77   n78 0      1f

R_78   n79 n78 1
C_78   n79 0      1f

R_79   n80 n79 1
C_79   n80 0      1f

R_80   n81 n80 1
C_80   n81 0      1f

R_81   n82 n81 1
C_81   n82 0      1f

R_82   n83 n82 1
C_82   n83 0      1f

R_83   n84 n83 1
C_83   n84 0      1f

R_84   n85 n84 1
C_84   n85 0      1f

R_85   n86 n85 1
C_85   n86 0      1f

R_86   n87 n86 1
C_86   n87 0      1f

R_87   n88 n87 1
C_87   n88 0      1f

R_88   n89 n88 1
C_88   n89 0      1f

R_89   n90 n89 1
C_89   n90 0      1f

R_90   n91 n90 1
C_90   n91 0      1f

R_91   n92 n91 1
C_91   n92 0      1f

R_92   n93 n92 1
C_92   n93 0      1f

R_93   n94 n93 1
C_93   n94 0      1f

R_94   n95 n94 1
C_94   n95 0      1f

R_95   n96 n95 1
C_95   n96 0      1f

R_96   n97 n96 1
C_96   n97 0      1f

R_97   n98 n97 1
C_97   n98 0      1f

R_98   n99 n98 1
C_98   n99 0      1f

R_99   n100 n99 1
C_99   n100 0      1f

R_100   n101 n100 1
C_100   n101 0      1f

R_101   n102 n101 1
C_101   n102 0      1f

R_102   n103 n102 1
C_102   n103 0      1f

R_103   n104 n103 1
C_103   n104 0      1f

R_104   n105 n104 1
C_104   n105 0      1f

R_105   n106 n105 1
C_105   n106 0      1f

R_106   n107 n106 1
C_106   n107 0      1f

R_107   n108 n107 1
C_107   n108 0      1f

R_108   n109 n108 1
C_108   n109 0      1f

R_109   n110 n109 1
C_109   n110 0      1f

R_110   n111 n110 1
C_110   n111 0      1f

R_111   n112 n111 1
C_111   n112 0      1f

R_112   n113 n112 1
C_112   n113 0      1f

R_113   n114 n113 1
C_113   n114 0      1f

R_114   n115 n114 1
C_114   n115 0      1f

R_115   n116 n115 1
C_115   n116 0      1f

R_116   n117 n116 1
C_116   n117 0      1f

R_117   n118 n117 1
C_117   n118 0      1f

R_118   n119 n118 1
C_118   n119 0      1f

R_119   n120 n119 1
C_119   n120 0      1f

R_120   n121 n120 1
C_120   n121 0      1f

R_121   n122 n121 1
C_121   n122 0      1f

R_122   n123 n122 1
C_122   n123 0      1f

R_123   n124 n123 1
C_123   n124 0      1f

R_124   n125 n124 1
C_124   n125 0      1f

R_125   n126 n125 1
C_125   n126 0      1f

R_126   n127 n126 1
C_126   n127 0      1f

R_127   n128 n127 1
C_127   n128 0      1f

R_128   n129 n128 1
C_128   n129 0      1f

R_129   n130 n129 1
C_129   n130 0      1f

R_130   n131 n130 1
C_130   n131 0      1f

R_131   n132 n131 1
C_131   n132 0      1f

R_132   n133 n132 1
C_132   n133 0      1f

R_133   n134 n133 1
C_133   n134 0      1f

R_134   n135 n134 1
C_134   n135 0      1f

R_135   n136 n135 1
C_135   n136 0      1f

R_136   n137 n136 1
C_136   n137 0      1f

R_137   n138 n137 1
C_137   n138 0      1f

R_138   n139 n138 1
C_138   n139 0      1f

R_139   n140 n139 1
C_139   n140 0      1f

R_140   n141 n140 1
C_140   n141 0      1f

R_141   n142 n141 1
C_141   n142 0      1f

R_142   n143 n142 1
C_142   n143 0      1f

R_143   n144 n143 1
C_143   n144 0      1f

R_144   n145 n144 1
C_144   n145 0      1f

R_145   n146 n145 1
C_145   n146 0      1f

R_146   n147 n146 1
C_146   n147 0      1f

R_147   n148 n147 1
C_147   n148 0      1f

R_148   n149 n148 1
C_148   n149 0      1f

R_149   n150 n149 1
C_149   n150 0      1f

R_150   n151 n150 1
C_150   n151 0      1f

R_151   n152 n151 1
C_151   n152 0      1f

R_152   n153 n152 1
C_152   n153 0      1f

R_153   n154 n153 1
C_153   n154 0      1f

R_154   n155 n154 1
C_154   n155 0      1f

R_155   n156 n155 1
C_155   n156 0      1f

R_156   n157 n156 1
C_156   n157 0      1f

R_157   n158 n157 1
C_157   n158 0      1f

R_158   n159 n158 1
C_158   n159 0      1f

R_159   n160 n159 1
C_159   n160 0      1f

R_160   n161 n160 1
C_160   n161 0      1f

R_161   n162 n161 1
C_161   n162 0      1f

R_162   n163 n162 1
C_162   n163 0      1f

R_163   n164 n163 1
C_163   n164 0      1f

R_164   n165 n164 1
C_164   n165 0      1f

R_165   n166 n165 1
C_165   n166 0      1f

R_166   n167 n166 1
C_166   n167 0      1f

R_167   n168 n167 1
C_167   n168 0      1f

R_168   n169 n168 1
C_168   n169 0      1f

R_169   n170 n169 1
C_169   n170 0      1f

R_170   n171 n170 1
C_170   n171 0      1f

R_171   n172 n171 1
C_171   n172 0      1f

R_172   n173 n172 1
C_172   n173 0      1f

R_173   n174 n173 1
C_173   n174 0      1f

R_174   n175 n174 1
C_174   n175 0      1f

R_175   n176 n175 1
C_175   n176 0      1f

R_176   n177 n176 1
C_176   n177 0      1f

R_177   n178 n177 1
C_177   n178 0      1f

R_178   n179 n178 1
C_178   n179 0      1f

R_179   n180 n179 1
C_179   n180 0      1f

R_180   n181 n180 1
C_180   n181 0      1f

R_181   n182 n181 1
C_181   n182 0      1f

R_182   n183 n182 1
C_182   n183 0      1f

R_183   n184 n183 1
C_183   n184 0      1f

R_184   n185 n184 1
C_184   n185 0      1f

R_185   n186 n185 1
C_185   n186 0      1f

R_186   n187 n186 1
C_186   n187 0      1f

R_187   n188 n187 1
C_187   n188 0      1f

R_188   n189 n188 1
C_188   n189 0      1f

R_189   n190 n189 1
C_189   n190 0      1f

R_190   n191 n190 1
C_190   n191 0      1f

R_191   n192 n191 1
C_191   n192 0      1f

R_192   n193 n192 1
C_192   n193 0      1f

R_193   n194 n193 1
C_193   n194 0      1f

R_194   n195 n194 1
C_194   n195 0      1f

R_195   n196 n195 1
C_195   n196 0      1f

R_196   n197 n196 1
C_196   n197 0      1f

R_197   n198 n197 1
C_197   n198 0      1f

R_198   n199 n198 1
C_198   n199 0      1f

R_199   n200 n199 1
C_199   n200 0      1f

R_200   n201 n200 1
C_200   n201 0      1f

R_201   n202 n201 1
C_201   n202 0      1f

R_202   n203 n202 1
C_202   n203 0      1f

R_203   n204 n203 1
C_203   n204 0      1f

R_204   n205 n204 1
C_204   n205 0      1f

R_205   n206 n205 1
C_205   n206 0      1f

R_206   n207 n206 1
C_206   n207 0      1f

R_207   n208 n207 1
C_207   n208 0      1f

R_208   n209 n208 1
C_208   n209 0      1f

R_209   n210 n209 1
C_209   n210 0      1f

R_210   n211 n210 1
C_210   n211 0      1f

R_211   n212 n211 1
C_211   n212 0      1f

R_212   n213 n212 1
C_212   n213 0      1f

R_213   n214 n213 1
C_213   n214 0      1f

R_214   n215 n214 1
C_214   n215 0      1f

R_215   n216 n215 1
C_215   n216 0      1f

R_216   n217 n216 1
C_216   n217 0      1f

R_217   n218 n217 1
C_217   n218 0      1f

R_218   n219 n218 1
C_218   n219 0      1f

R_219   n220 n219 1
C_219   n220 0      1f

R_220   n221 n220 1
C_220   n221 0      1f

R_221   n222 n221 1
C_221   n222 0      1f

R_222   n223 n222 1
C_222   n223 0      1f

R_223   n224 n223 1
C_223   n224 0      1f

R_224   n225 n224 1
C_224   n225 0      1f

R_225   n226 n225 1
C_225   n226 0      1f

R_226   n227 n226 1
C_226   n227 0      1f

R_227   n228 n227 1
C_227   n228 0      1f

R_228   n229 n228 1
C_228   n229 0      1f

R_229   n230 n229 1
C_229   n230 0      1f

R_230   n231 n230 1
C_230   n231 0      1f

R_231   n232 n231 1
C_231   n232 0      1f

R_232   n233 n232 1
C_232   n233 0      1f

R_233   n234 n233 1
C_233   n234 0      1f

R_234   n235 n234 1
C_234   n235 0      1f

R_235   n236 n235 1
C_235   n236 0      1f

R_236   n237 n236 1
C_236   n237 0      1f

R_237   n238 n237 1
C_237   n238 0      1f

R_238   n239 n238 1
C_238   n239 0      1f

R_239   n240 n239 1
C_239   n240 0      1f

R_240   n241 n240 1
C_240   n241 0      1f

R_241   n242 n241 1
C_241   n242 0      1f

R_242   n243 n242 1
C_242   n243 0      1f

R_243   n244 n243 1
C_243   n244 0      1f

R_244   n245 n244 1
C_244   n245 0      1f

R_245   n246 n245 1
C_245   n246 0      1f

R_246   n247 n246 1
C_246   n247 0      1f

R_247   n248 n247 1
C_247   n248 0      1f

R_248   n249 n248 1
C_248   n249 0      1f

R_249   n250 n249 1
C_249   n250 0      1f

R_250   n251 n250 1
C_250   n251 0      1f

R_251   n252 n251 1
C_251   n252 0      1f

R_252   n253 n252 1
C_252   n253 0      1f

R_253   n254 n253 1
C_253   n254 0      1f

R_254   n255 n254 1
C_254   n255 0      1f

R_255   n256 n255 1
C_255   n256 0      1f

R_256   n257 n256 1
C_256   n257 0      1f

R_257   n258 n257 1
C_257   n258 0      1f

R_258   n259 n258 1
C_258   n259 0      1f

R_259   n260 n259 1
C_259   n260 0      1f

R_260   n261 n260 1
C_260   n261 0      1f

R_261   n262 n261 1
C_261   n262 0      1f

R_262   n263 n262 1
C_262   n263 0      1f

R_263   n264 n263 1
C_263   n264 0      1f

R_264   n265 n264 1
C_264   n265 0      1f

R_265   n266 n265 1
C_265   n266 0      1f

R_266   n267 n266 1
C_266   n267 0      1f

R_267   n268 n267 1
C_267   n268 0      1f

R_268   n269 n268 1
C_268   n269 0      1f

R_269   n270 n269 1
C_269   n270 0      1f

R_270   n271 n270 1
C_270   n271 0      1f

R_271   n272 n271 1
C_271   n272 0      1f

R_272   n273 n272 1
C_272   n273 0      1f

R_273   n274 n273 1
C_273   n274 0      1f

R_274   n275 n274 1
C_274   n275 0      1f

R_275   n276 n275 1
C_275   n276 0      1f

R_276   n277 n276 1
C_276   n277 0      1f

R_277   n278 n277 1
C_277   n278 0      1f

R_278   n279 n278 1
C_278   n279 0      1f

R_279   n280 n279 1
C_279   n280 0      1f

R_280   n281 n280 1
C_280   n281 0      1f

R_281   n282 n281 1
C_281   n282 0      1f

R_282   n283 n282 1
C_282   n283 0      1f

R_283   n284 n283 1
C_283   n284 0      1f

R_284   n285 n284 1
C_284   n285 0      1f

R_285   n286 n285 1
C_285   n286 0      1f

R_286   n287 n286 1
C_286   n287 0      1f

R_287   n288 n287 1
C_287   n288 0      1f

R_288   n289 n288 1
C_288   n289 0      1f

R_289   n290 n289 1
C_289   n290 0      1f

R_290   n291 n290 1
C_290   n291 0      1f

R_291   n292 n291 1
C_291   n292 0      1f

R_292   n293 n292 1
C_292   n293 0      1f

R_293   n294 n293 1
C_293   n294 0      1f

R_294   n295 n294 1
C_294   n295 0      1f

R_295   n296 n295 1
C_295   n296 0      1f

R_296   n297 n296 1
C_296   n297 0      1f

R_297   n298 n297 1
C_297   n298 0      1f

R_298   n299 n298 1
C_298   n299 0      1f

R_299   n300 n299 1
C_299   n300 0      1f

R_300   n301 n300 1
C_300   n301 0      1f

R_301   n302 n301 1
C_301   n302 0      1f

R_302   n303 n302 1
C_302   n303 0      1f

R_303   n304 n303 1
C_303   n304 0      1f

R_304   n305 n304 1
C_304   n305 0      1f

R_305   n306 n305 1
C_305   n306 0      1f

R_306   n307 n306 1
C_306   n307 0      1f

R_307   n308 n307 1
C_307   n308 0      1f

R_308   n309 n308 1
C_308   n309 0      1f

R_309   n310 n309 1
C_309   n310 0      1f

R_310   n311 n310 1
C_310   n311 0      1f

R_311   n312 n311 1
C_311   n312 0      1f

R_312   n313 n312 1
C_312   n313 0      1f

R_313   n314 n313 1
C_313   n314 0      1f

R_314   n315 n314 1
C_314   n315 0      1f

R_315   n316 n315 1
C_315   n316 0      1f

R_316   n317 n316 1
C_316   n317 0      1f

R_317   n318 n317 1
C_317   n318 0      1f

R_318   n319 n318 1
C_318   n319 0      1f

R_319   n320 n319 1
C_319   n320 0      1f

R_320   n321 n320 1
C_320   n321 0      1f

R_321   n322 n321 1
C_321   n322 0      1f

R_322   n323 n322 1
C_322   n323 0      1f

R_323   n324 n323 1
C_323   n324 0      1f

R_324   n325 n324 1
C_324   n325 0      1f

R_325   n326 n325 1
C_325   n326 0      1f

R_326   n327 n326 1
C_326   n327 0      1f

R_327   n328 n327 1
C_327   n328 0      1f

R_328   n329 n328 1
C_328   n329 0      1f

R_329   n330 n329 1
C_329   n330 0      1f

R_330   n331 n330 1
C_330   n331 0      1f

R_331   n332 n331 1
C_331   n332 0      1f

R_332   n333 n332 1
C_332   n333 0      1f

R_333   n334 n333 1
C_333   n334 0      1f

R_334   n335 n334 1
C_334   n335 0      1f

R_335   n336 n335 1
C_335   n336 0      1f

R_336   n337 n336 1
C_336   n337 0      1f

R_337   n338 n337 1
C_337   n338 0      1f

R_338   n339 n338 1
C_338   n339 0      1f

R_339   n340 n339 1
C_339   n340 0      1f

R_340   n341 n340 1
C_340   n341 0      1f

R_341   n342 n341 1
C_341   n342 0      1f

R_342   n343 n342 1
C_342   n343 0      1f

R_343   n344 n343 1
C_343   n344 0      1f

R_344   n345 n344 1
C_344   n345 0      1f

R_345   n346 n345 1
C_345   n346 0      1f

R_346   n347 n346 1
C_346   n347 0      1f

R_347   n348 n347 1
C_347   n348 0      1f

R_348   n349 n348 1
C_348   n349 0      1f

R_349   n350 n349 1
C_349   n350 0      1f

R_350   n351 n350 1
C_350   n351 0      1f

R_351   n352 n351 1
C_351   n352 0      1f

R_352   n353 n352 1
C_352   n353 0      1f

R_353   n354 n353 1
C_353   n354 0      1f

R_354   n355 n354 1
C_354   n355 0      1f

R_355   n356 n355 1
C_355   n356 0      1f

R_356   n357 n356 1
C_356   n357 0      1f

R_357   n358 n357 1
C_357   n358 0      1f

R_358   n359 n358 1
C_358   n359 0      1f

R_359   n360 n359 1
C_359   n360 0      1f

R_360   n361 n360 1
C_360   n361 0      1f

R_361   n362 n361 1
C_361   n362 0      1f

R_362   n363 n362 1
C_362   n363 0      1f

R_363   n364 n363 1
C_363   n364 0      1f

R_364   n365 n364 1
C_364   n365 0      1f

R_365   n366 n365 1
C_365   n366 0      1f

R_366   n367 n366 1
C_366   n367 0      1f

R_367   n368 n367 1
C_367   n368 0      1f

R_368   n369 n368 1
C_368   n369 0      1f

R_369   n370 n369 1
C_369   n370 0      1f

R_370   n371 n370 1
C_370   n371 0      1f

R_371   n372 n371 1
C_371   n372 0      1f

R_372   n373 n372 1
C_372   n373 0      1f

R_373   n374 n373 1
C_373   n374 0      1f

R_374   n375 n374 1
C_374   n375 0      1f

R_375   n376 n375 1
C_375   n376 0      1f

R_376   n377 n376 1
C_376   n377 0      1f

R_377   n378 n377 1
C_377   n378 0      1f

R_378   n379 n378 1
C_378   n379 0      1f

R_379   n380 n379 1
C_379   n380 0      1f

R_380   n381 n380 1
C_380   n381 0      1f

R_381   n382 n381 1
C_381   n382 0      1f

R_382   n383 n382 1
C_382   n383 0      1f

R_383   n384 n383 1
C_383   n384 0      1f

R_384   n385 n384 1
C_384   n385 0      1f

R_385   n386 n385 1
C_385   n386 0      1f

R_386   n387 n386 1
C_386   n387 0      1f

R_387   n388 n387 1
C_387   n388 0      1f

R_388   n389 n388 1
C_388   n389 0      1f

R_389   n390 n389 1
C_389   n390 0      1f

R_390   n391 n390 1
C_390   n391 0      1f

R_391   n392 n391 1
C_391   n392 0      1f

R_392   n393 n392 1
C_392   n393 0      1f

R_393   n394 n393 1
C_393   n394 0      1f

R_394   n395 n394 1
C_394   n395 0      1f

R_395   n396 n395 1
C_395   n396 0      1f

R_396   n397 n396 1
C_396   n397 0      1f

R_397   n398 n397 1
C_397   n398 0      1f

R_398   n399 n398 1
C_398   n399 0      1f

R_399   n400 n399 1
C_399   n400 0      1f

R_400   n401 n400 1
C_400   n401 0      1f

R_401   n402 n401 1
C_401   n402 0      1f

R_402   n403 n402 1
C_402   n403 0      1f

R_403   n404 n403 1
C_403   n404 0      1f

R_404   n405 n404 1
C_404   n405 0      1f

R_405   n406 n405 1
C_405   n406 0      1f

R_406   n407 n406 1
C_406   n407 0      1f

R_407   n408 n407 1
C_407   n408 0      1f

R_408   n409 n408 1
C_408   n409 0      1f

R_409   n410 n409 1
C_409   n410 0      1f

R_410   n411 n410 1
C_410   n411 0      1f

R_411   n412 n411 1
C_411   n412 0      1f

R_412   n413 n412 1
C_412   n413 0      1f

R_413   n414 n413 1
C_413   n414 0      1f

R_414   n415 n414 1
C_414   n415 0      1f

R_415   n416 n415 1
C_415   n416 0      1f

R_416   n417 n416 1
C_416   n417 0      1f

R_417   n418 n417 1
C_417   n418 0      1f

R_418   n419 n418 1
C_418   n419 0      1f

R_419   n420 n419 1
C_419   n420 0      1f

R_420   n421 n420 1
C_420   n421 0      1f

R_421   n422 n421 1
C_421   n422 0      1f

R_422   n423 n422 1
C_422   n423 0      1f

R_423   n424 n423 1
C_423   n424 0      1f

R_424   n425 n424 1
C_424   n425 0      1f

R_425   n426 n425 1
C_425   n426 0      1f

R_426   n427 n426 1
C_426   n427 0      1f

R_427   n428 n427 1
C_427   n428 0      1f

R_428   n429 n428 1
C_428   n429 0      1f

R_429   n430 n429 1
C_429   n430 0      1f

R_430   n431 n430 1
C_430   n431 0      1f

R_431   n432 n431 1
C_431   n432 0      1f

R_432   n433 n432 1
C_432   n433 0      1f

R_433   n434 n433 1
C_433   n434 0      1f

R_434   n435 n434 1
C_434   n435 0      1f

R_435   n436 n435 1
C_435   n436 0      1f

R_436   n437 n436 1
C_436   n437 0      1f

R_437   n438 n437 1
C_437   n438 0      1f

R_438   n439 n438 1
C_438   n439 0      1f

R_439   n440 n439 1
C_439   n440 0      1f

R_440   n441 n440 1
C_440   n441 0      1f

R_441   n442 n441 1
C_441   n442 0      1f

R_442   n443 n442 1
C_442   n443 0      1f

R_443   n444 n443 1
C_443   n444 0      1f

R_444   n445 n444 1
C_444   n445 0      1f

R_445   n446 n445 1
C_445   n446 0      1f

R_446   n447 n446 1
C_446   n447 0      1f

R_447   n448 n447 1
C_447   n448 0      1f

R_448   n449 n448 1
C_448   n449 0      1f

R_449   n450 n449 1
C_449   n450 0      1f

R_450   n451 n450 1
C_450   n451 0      1f

R_451   n452 n451 1
C_451   n452 0      1f

R_452   n453 n452 1
C_452   n453 0      1f

R_453   n454 n453 1
C_453   n454 0      1f

R_454   n455 n454 1
C_454   n455 0      1f

R_455   n456 n455 1
C_455   n456 0      1f

R_456   n457 n456 1
C_456   n457 0      1f

R_457   n458 n457 1
C_457   n458 0      1f

R_458   n459 n458 1
C_458   n459 0      1f

R_459   n460 n459 1
C_459   n460 0      1f

R_460   n461 n460 1
C_460   n461 0      1f

R_461   n462 n461 1
C_461   n462 0      1f

R_462   n463 n462 1
C_462   n463 0      1f

R_463   n464 n463 1
C_463   n464 0      1f

R_464   n465 n464 1
C_464   n465 0      1f

R_465   n466 n465 1
C_465   n466 0      1f

R_466   n467 n466 1
C_466   n467 0      1f

R_467   n468 n467 1
C_467   n468 0      1f

R_468   n469 n468 1
C_468   n469 0      1f

R_469   n470 n469 1
C_469   n470 0      1f

R_470   n471 n470 1
C_470   n471 0      1f

R_471   n472 n471 1
C_471   n472 0      1f

R_472   n473 n472 1
C_472   n473 0      1f

R_473   n474 n473 1
C_473   n474 0      1f

R_474   n475 n474 1
C_474   n475 0      1f

R_475   n476 n475 1
C_475   n476 0      1f

R_476   n477 n476 1
C_476   n477 0      1f

R_477   n478 n477 1
C_477   n478 0      1f

R_478   n479 n478 1
C_478   n479 0      1f

R_479   n480 n479 1
C_479   n480 0      1f

R_480   n481 n480 1
C_480   n481 0      1f

R_481   n482 n481 1
C_481   n482 0      1f

R_482   n483 n482 1
C_482   n483 0      1f

R_483   n484 n483 1
C_483   n484 0      1f

R_484   n485 n484 1
C_484   n485 0      1f

R_485   n486 n485 1
C_485   n486 0      1f

R_486   n487 n486 1
C_486   n487 0      1f

R_487   n488 n487 1
C_487   n488 0      1f

R_488   n489 n488 1
C_488   n489 0      1f

R_489   n490 n489 1
C_489   n490 0      1f

R_490   n491 n490 1
C_490   n491 0      1f

R_491   n492 n491 1
C_491   n492 0      1f

R_492   n493 n492 1
C_492   n493 0      1f

R_493   n494 n493 1
C_493   n494 0      1f

R_494   n495 n494 1
C_494   n495 0      1f

R_495   n496 n495 1
C_495   n496 0      1f

R_496   n497 n496 1
C_496   n497 0      1f

R_497   n498 n497 1
C_497   n498 0      1f

R_498   n499 n498 1
C_498   n499 0      1f

R_499   n500 n499 1
C_499   n500 0      1f

R_500   n501 n500 1
C_500   n501 0      1f

R_501   n502 n501 1
C_501   n502 0      1f

R_502   n503 n502 1
C_502   n503 0      1f

R_503   n504 n503 1
C_503   n504 0      1f

R_504   n505 n504 1
C_504   n505 0      1f

R_505   n506 n505 1
C_505   n506 0      1f

R_506   n507 n506 1
C_506   n507 0      1f

R_507   n508 n507 1
C_507   n508 0      1f

R_508   n509 n508 1
C_508   n509 0      1f

R_509   n510 n509 1
C_509   n510 0      1f

R_510   n511 n510 1
C_510   n511 0      1f

R_511   n512 n511 1
C_511   n512 0      1f

R_512   n513 n512 1
C_512   n513 0      1f

R_513   n514 n513 1
C_513   n514 0      1f

R_514   n515 n514 1
C_514   n515 0      1f

R_515   n516 n515 1
C_515   n516 0      1f

R_516   n517 n516 1
C_516   n517 0      1f

R_517   n518 n517 1
C_517   n518 0      1f

R_518   n519 n518 1
C_518   n519 0      1f

R_519   n520 n519 1
C_519   n520 0      1f

R_520   n521 n520 1
C_520   n521 0      1f

R_521   n522 n521 1
C_521   n522 0      1f

R_522   n523 n522 1
C_522   n523 0      1f

R_523   n524 n523 1
C_523   n524 0      1f

R_524   n525 n524 1
C_524   n525 0      1f

R_525   n526 n525 1
C_525   n526 0      1f

R_526   n527 n526 1
C_526   n527 0      1f

R_527   n528 n527 1
C_527   n528 0      1f

R_528   n529 n528 1
C_528   n529 0      1f

R_529   n530 n529 1
C_529   n530 0      1f

R_530   n531 n530 1
C_530   n531 0      1f

R_531   n532 n531 1
C_531   n532 0      1f

R_532   n533 n532 1
C_532   n533 0      1f

R_533   n534 n533 1
C_533   n534 0      1f

R_534   n535 n534 1
C_534   n535 0      1f

R_535   n536 n535 1
C_535   n536 0      1f

R_536   n537 n536 1
C_536   n537 0      1f

R_537   n538 n537 1
C_537   n538 0      1f

R_538   n539 n538 1
C_538   n539 0      1f

R_539   n540 n539 1
C_539   n540 0      1f

R_540   n541 n540 1
C_540   n541 0      1f

R_541   n542 n541 1
C_541   n542 0      1f

R_542   n543 n542 1
C_542   n543 0      1f

R_543   n544 n543 1
C_543   n544 0      1f

R_544   n545 n544 1
C_544   n545 0      1f

R_545   n546 n545 1
C_545   n546 0      1f

R_546   n547 n546 1
C_546   n547 0      1f

R_547   n548 n547 1
C_547   n548 0      1f

R_548   n549 n548 1
C_548   n549 0      1f

R_549   n550 n549 1
C_549   n550 0      1f

R_550   n551 n550 1
C_550   n551 0      1f

R_551   n552 n551 1
C_551   n552 0      1f

R_552   n553 n552 1
C_552   n553 0      1f

R_553   n554 n553 1
C_553   n554 0      1f

R_554   n555 n554 1
C_554   n555 0      1f

R_555   n556 n555 1
C_555   n556 0      1f

R_556   n557 n556 1
C_556   n557 0      1f

R_557   n558 n557 1
C_557   n558 0      1f

R_558   n559 n558 1
C_558   n559 0      1f

R_559   n560 n559 1
C_559   n560 0      1f

R_560   n561 n560 1
C_560   n561 0      1f

R_561   n562 n561 1
C_561   n562 0      1f

R_562   n563 n562 1
C_562   n563 0      1f

R_563   n564 n563 1
C_563   n564 0      1f

R_564   n565 n564 1
C_564   n565 0      1f

R_565   n566 n565 1
C_565   n566 0      1f

R_566   n567 n566 1
C_566   n567 0      1f

R_567   n568 n567 1
C_567   n568 0      1f

R_568   n569 n568 1
C_568   n569 0      1f

R_569   n570 n569 1
C_569   n570 0      1f

R_570   n571 n570 1
C_570   n571 0      1f

R_571   n572 n571 1
C_571   n572 0      1f

R_572   n573 n572 1
C_572   n573 0      1f

R_573   n574 n573 1
C_573   n574 0      1f

R_574   n575 n574 1
C_574   n575 0      1f

R_575   n576 n575 1
C_575   n576 0      1f

R_576   n577 n576 1
C_576   n577 0      1f

R_577   n578 n577 1
C_577   n578 0      1f

R_578   n579 n578 1
C_578   n579 0      1f

R_579   n580 n579 1
C_579   n580 0      1f

R_580   n581 n580 1
C_580   n581 0      1f

R_581   n582 n581 1
C_581   n582 0      1f

R_582   n583 n582 1
C_582   n583 0      1f

R_583   n584 n583 1
C_583   n584 0      1f

R_584   n585 n584 1
C_584   n585 0      1f

R_585   n586 n585 1
C_585   n586 0      1f

R_586   n587 n586 1
C_586   n587 0      1f

R_587   n588 n587 1
C_587   n588 0      1f

R_588   n589 n588 1
C_588   n589 0      1f

R_589   n590 n589 1
C_589   n590 0      1f

R_590   n591 n590 1
C_590   n591 0      1f

R_591   n592 n591 1
C_591   n592 0      1f

R_592   n593 n592 1
C_592   n593 0      1f

R_593   n594 n593 1
C_593   n594 0      1f

R_594   n595 n594 1
C_594   n595 0      1f

R_595   n596 n595 1
C_595   n596 0      1f

R_596   n597 n596 1
C_596   n597 0      1f

R_597   n598 n597 1
C_597   n598 0      1f

R_598   n599 n598 1
C_598   n599 0      1f

R_599   n600 n599 1
C_599   n600 0      1f

R_600   n601 n600 1
C_600   n601 0      1f

R_601   n602 n601 1
C_601   n602 0      1f

R_602   n603 n602 1
C_602   n603 0      1f

R_603   n604 n603 1
C_603   n604 0      1f

R_604   n605 n604 1
C_604   n605 0      1f

R_605   n606 n605 1
C_605   n606 0      1f

R_606   n607 n606 1
C_606   n607 0      1f

R_607   n608 n607 1
C_607   n608 0      1f

R_608   n609 n608 1
C_608   n609 0      1f

R_609   n610 n609 1
C_609   n610 0      1f

R_610   n611 n610 1
C_610   n611 0      1f

R_611   n612 n611 1
C_611   n612 0      1f

R_612   n613 n612 1
C_612   n613 0      1f

R_613   n614 n613 1
C_613   n614 0      1f

R_614   n615 n614 1
C_614   n615 0      1f

R_615   n616 n615 1
C_615   n616 0      1f

R_616   n617 n616 1
C_616   n617 0      1f

R_617   n618 n617 1
C_617   n618 0      1f

R_618   n619 n618 1
C_618   n619 0      1f

R_619   n620 n619 1
C_619   n620 0      1f

R_620   n621 n620 1
C_620   n621 0      1f

R_621   n622 n621 1
C_621   n622 0      1f

R_622   n623 n622 1
C_622   n623 0      1f

R_623   n624 n623 1
C_623   n624 0      1f

R_624   n625 n624 1
C_624   n625 0      1f

R_625   n626 n625 1
C_625   n626 0      1f

R_626   n627 n626 1
C_626   n627 0      1f

R_627   n628 n627 1
C_627   n628 0      1f

R_628   n629 n628 1
C_628   n629 0      1f

R_629   n630 n629 1
C_629   n630 0      1f

R_630   n631 n630 1
C_630   n631 0      1f

R_631   n632 n631 1
C_631   n632 0      1f

R_632   n633 n632 1
C_632   n633 0      1f

R_633   n634 n633 1
C_633   n634 0      1f

R_634   n635 n634 1
C_634   n635 0      1f

R_635   n636 n635 1
C_635   n636 0      1f

R_636   n637 n636 1
C_636   n637 0      1f

R_637   n638 n637 1
C_637   n638 0      1f

R_638   n639 n638 1
C_638   n639 0      1f

R_639   n640 n639 1
C_639   n640 0      1f

R_640   n641 n640 1
C_640   n641 0      1f

R_641   n642 n641 1
C_641   n642 0      1f

R_642   n643 n642 1
C_642   n643 0      1f

R_643   n644 n643 1
C_643   n644 0      1f

R_644   n645 n644 1
C_644   n645 0      1f

R_645   n646 n645 1
C_645   n646 0      1f

R_646   n647 n646 1
C_646   n647 0      1f

R_647   n648 n647 1
C_647   n648 0      1f

R_648   n649 n648 1
C_648   n649 0      1f

R_649   n650 n649 1
C_649   n650 0      1f

R_650   n651 n650 1
C_650   n651 0      1f

R_651   n652 n651 1
C_651   n652 0      1f

R_652   n653 n652 1
C_652   n653 0      1f

R_653   n654 n653 1
C_653   n654 0      1f

R_654   n655 n654 1
C_654   n655 0      1f

R_655   n656 n655 1
C_655   n656 0      1f

R_656   n657 n656 1
C_656   n657 0      1f

R_657   n658 n657 1
C_657   n658 0      1f

R_658   n659 n658 1
C_658   n659 0      1f

R_659   n660 n659 1
C_659   n660 0      1f

R_660   n661 n660 1
C_660   n661 0      1f

R_661   n662 n661 1
C_661   n662 0      1f

R_662   n663 n662 1
C_662   n663 0      1f

R_663   n664 n663 1
C_663   n664 0      1f

R_664   n665 n664 1
C_664   n665 0      1f

R_665   n666 n665 1
C_665   n666 0      1f

R_666   n667 n666 1
C_666   n667 0      1f

R_667   n668 n667 1
C_667   n668 0      1f

R_668   n669 n668 1
C_668   n669 0      1f

R_669   n670 n669 1
C_669   n670 0      1f

R_670   n671 n670 1
C_670   n671 0      1f

R_671   n672 n671 1
C_671   n672 0      1f

R_672   n673 n672 1
C_672   n673 0      1f

R_673   n674 n673 1
C_673   n674 0      1f

R_674   n675 n674 1
C_674   n675 0      1f

R_675   n676 n675 1
C_675   n676 0      1f

R_676   n677 n676 1
C_676   n677 0      1f

R_677   n678 n677 1
C_677   n678 0      1f

R_678   n679 n678 1
C_678   n679 0      1f

R_679   n680 n679 1
C_679   n680 0      1f

R_680   n681 n680 1
C_680   n681 0      1f

R_681   n682 n681 1
C_681   n682 0      1f

R_682   n683 n682 1
C_682   n683 0      1f

R_683   n684 n683 1
C_683   n684 0      1f

R_684   n685 n684 1
C_684   n685 0      1f

R_685   n686 n685 1
C_685   n686 0      1f

R_686   n687 n686 1
C_686   n687 0      1f

R_687   n688 n687 1
C_687   n688 0      1f

R_688   n689 n688 1
C_688   n689 0      1f

R_689   n690 n689 1
C_689   n690 0      1f

R_690   n691 n690 1
C_690   n691 0      1f

R_691   n692 n691 1
C_691   n692 0      1f

R_692   n693 n692 1
C_692   n693 0      1f

R_693   n694 n693 1
C_693   n694 0      1f

R_694   n695 n694 1
C_694   n695 0      1f

R_695   n696 n695 1
C_695   n696 0      1f

R_696   n697 n696 1
C_696   n697 0      1f

R_697   n698 n697 1
C_697   n698 0      1f

R_698   n699 n698 1
C_698   n699 0      1f

R_699   n700 n699 1
C_699   n700 0      1f

R_700   n701 n700 1
C_700   n701 0      1f

R_701   n702 n701 1
C_701   n702 0      1f

R_702   n703 n702 1
C_702   n703 0      1f

R_703   n704 n703 1
C_703   n704 0      1f

R_704   n705 n704 1
C_704   n705 0      1f

R_705   n706 n705 1
C_705   n706 0      1f

R_706   n707 n706 1
C_706   n707 0      1f

R_707   n708 n707 1
C_707   n708 0      1f

R_708   n709 n708 1
C_708   n709 0      1f

R_709   n710 n709 1
C_709   n710 0      1f

R_710   n711 n710 1
C_710   n711 0      1f

R_711   n712 n711 1
C_711   n712 0      1f

R_712   n713 n712 1
C_712   n713 0      1f

R_713   n714 n713 1
C_713   n714 0      1f

R_714   n715 n714 1
C_714   n715 0      1f

R_715   n716 n715 1
C_715   n716 0      1f

R_716   n717 n716 1
C_716   n717 0      1f

R_717   n718 n717 1
C_717   n718 0      1f

R_718   n719 n718 1
C_718   n719 0      1f

R_719   n720 n719 1
C_719   n720 0      1f

R_720   n721 n720 1
C_720   n721 0      1f

R_721   n722 n721 1
C_721   n722 0      1f

R_722   n723 n722 1
C_722   n723 0      1f

R_723   n724 n723 1
C_723   n724 0      1f

R_724   n725 n724 1
C_724   n725 0      1f

R_725   n726 n725 1
C_725   n726 0      1f

R_726   n727 n726 1
C_726   n727 0      1f

R_727   n728 n727 1
C_727   n728 0      1f

R_728   n729 n728 1
C_728   n729 0      1f

R_729   n730 n729 1
C_729   n730 0      1f

R_730   n731 n730 1
C_730   n731 0      1f

R_731   n732 n731 1
C_731   n732 0      1f

R_732   n733 n732 1
C_732   n733 0      1f

R_733   n734 n733 1
C_733   n734 0      1f

R_734   n735 n734 1
C_734   n735 0      1f

R_735   n736 n735 1
C_735   n736 0      1f

R_736   n737 n736 1
C_736   n737 0      1f

R_737   n738 n737 1
C_737   n738 0      1f

R_738   n739 n738 1
C_738   n739 0      1f

R_739   n740 n739 1
C_739   n740 0      1f

R_740   n741 n740 1
C_740   n741 0      1f

R_741   n742 n741 1
C_741   n742 0      1f

R_742   n743 n742 1
C_742   n743 0      1f

R_743   n744 n743 1
C_743   n744 0      1f

R_744   n745 n744 1
C_744   n745 0      1f

R_745   n746 n745 1
C_745   n746 0      1f

R_746   n747 n746 1
C_746   n747 0      1f

R_747   n748 n747 1
C_747   n748 0      1f

R_748   n749 n748 1
C_748   n749 0      1f

R_749   n750 n749 1
C_749   n750 0      1f

R_750   n751 n750 1
C_750   n751 0      1f

R_751   n752 n751 1
C_751   n752 0      1f

R_752   n753 n752 1
C_752   n753 0      1f

R_753   n754 n753 1
C_753   n754 0      1f

R_754   n755 n754 1
C_754   n755 0      1f

R_755   n756 n755 1
C_755   n756 0      1f

R_756   n757 n756 1
C_756   n757 0      1f

R_757   n758 n757 1
C_757   n758 0      1f

R_758   n759 n758 1
C_758   n759 0      1f

R_759   n760 n759 1
C_759   n760 0      1f

R_760   n761 n760 1
C_760   n761 0      1f

R_761   n762 n761 1
C_761   n762 0      1f

R_762   n763 n762 1
C_762   n763 0      1f

R_763   n764 n763 1
C_763   n764 0      1f

R_764   n765 n764 1
C_764   n765 0      1f

R_765   n766 n765 1
C_765   n766 0      1f

R_766   n767 n766 1
C_766   n767 0      1f

R_767   n768 n767 1
C_767   n768 0      1f

R_768   n769 n768 1
C_768   n769 0      1f

R_769   n770 n769 1
C_769   n770 0      1f

R_770   n771 n770 1
C_770   n771 0      1f

R_771   n772 n771 1
C_771   n772 0      1f

R_772   n773 n772 1
C_772   n773 0      1f

R_773   n774 n773 1
C_773   n774 0      1f

R_774   n775 n774 1
C_774   n775 0      1f

R_775   n776 n775 1
C_775   n776 0      1f

R_776   n777 n776 1
C_776   n777 0      1f

R_777   n778 n777 1
C_777   n778 0      1f

R_778   n779 n778 1
C_778   n779 0      1f

R_779   n780 n779 1
C_779   n780 0      1f

R_780   n781 n780 1
C_780   n781 0      1f

R_781   n782 n781 1
C_781   n782 0      1f

R_782   n783 n782 1
C_782   n783 0      1f

R_783   n784 n783 1
C_783   n784 0      1f

R_784   n785 n784 1
C_784   n785 0      1f

R_785   n786 n785 1
C_785   n786 0      1f

R_786   n787 n786 1
C_786   n787 0      1f

R_787   n788 n787 1
C_787   n788 0      1f

R_788   n789 n788 1
C_788   n789 0      1f

R_789   n790 n789 1
C_789   n790 0      1f

R_790   n791 n790 1
C_790   n791 0      1f

R_791   n792 n791 1
C_791   n792 0      1f

R_792   n793 n792 1
C_792   n793 0      1f

R_793   n794 n793 1
C_793   n794 0      1f

R_794   n795 n794 1
C_794   n795 0      1f

R_795   n796 n795 1
C_795   n796 0      1f

R_796   n797 n796 1
C_796   n797 0      1f

R_797   n798 n797 1
C_797   n798 0      1f

R_798   n799 n798 1
C_798   n799 0      1f

R_799   n800 n799 1
C_799   n800 0      1f

R_800   n801 n800 1
C_800   n801 0      1f

R_801   n802 n801 1
C_801   n802 0      1f

R_802   n803 n802 1
C_802   n803 0      1f

R_803   n804 n803 1
C_803   n804 0      1f

R_804   n805 n804 1
C_804   n805 0      1f

R_805   n806 n805 1
C_805   n806 0      1f

R_806   n807 n806 1
C_806   n807 0      1f

R_807   n808 n807 1
C_807   n808 0      1f

R_808   n809 n808 1
C_808   n809 0      1f

R_809   n810 n809 1
C_809   n810 0      1f

R_810   n811 n810 1
C_810   n811 0      1f

R_811   n812 n811 1
C_811   n812 0      1f

R_812   n813 n812 1
C_812   n813 0      1f

R_813   n814 n813 1
C_813   n814 0      1f

R_814   n815 n814 1
C_814   n815 0      1f

R_815   n816 n815 1
C_815   n816 0      1f

R_816   n817 n816 1
C_816   n817 0      1f

R_817   n818 n817 1
C_817   n818 0      1f

R_818   n819 n818 1
C_818   n819 0      1f

R_819   n820 n819 1
C_819   n820 0      1f

R_820   n821 n820 1
C_820   n821 0      1f

R_821   n822 n821 1
C_821   n822 0      1f

R_822   n823 n822 1
C_822   n823 0      1f

R_823   n824 n823 1
C_823   n824 0      1f

R_824   n825 n824 1
C_824   n825 0      1f

R_825   n826 n825 1
C_825   n826 0      1f

R_826   n827 n826 1
C_826   n827 0      1f

R_827   n828 n827 1
C_827   n828 0      1f

R_828   n829 n828 1
C_828   n829 0      1f

R_829   n830 n829 1
C_829   n830 0      1f

R_830   n831 n830 1
C_830   n831 0      1f

R_831   n832 n831 1
C_831   n832 0      1f

R_832   n833 n832 1
C_832   n833 0      1f

R_833   n834 n833 1
C_833   n834 0      1f

R_834   n835 n834 1
C_834   n835 0      1f

R_835   n836 n835 1
C_835   n836 0      1f

R_836   n837 n836 1
C_836   n837 0      1f

R_837   n838 n837 1
C_837   n838 0      1f

R_838   n839 n838 1
C_838   n839 0      1f

R_839   n840 n839 1
C_839   n840 0      1f

R_840   n841 n840 1
C_840   n841 0      1f

R_841   n842 n841 1
C_841   n842 0      1f

R_842   n843 n842 1
C_842   n843 0      1f

R_843   n844 n843 1
C_843   n844 0      1f

R_844   n845 n844 1
C_844   n845 0      1f

R_845   n846 n845 1
C_845   n846 0      1f

R_846   n847 n846 1
C_846   n847 0      1f

R_847   n848 n847 1
C_847   n848 0      1f

R_848   n849 n848 1
C_848   n849 0      1f

R_849   n850 n849 1
C_849   n850 0      1f

R_850   n851 n850 1
C_850   n851 0      1f

R_851   n852 n851 1
C_851   n852 0      1f

R_852   n853 n852 1
C_852   n853 0      1f

R_853   n854 n853 1
C_853   n854 0      1f

R_854   n855 n854 1
C_854   n855 0      1f

R_855   n856 n855 1
C_855   n856 0      1f

R_856   n857 n856 1
C_856   n857 0      1f

R_857   n858 n857 1
C_857   n858 0      1f

R_858   n859 n858 1
C_858   n859 0      1f

R_859   n860 n859 1
C_859   n860 0      1f

R_860   n861 n860 1
C_860   n861 0      1f

R_861   n862 n861 1
C_861   n862 0      1f

R_862   n863 n862 1
C_862   n863 0      1f

R_863   n864 n863 1
C_863   n864 0      1f

R_864   n865 n864 1
C_864   n865 0      1f

R_865   n866 n865 1
C_865   n866 0      1f

R_866   n867 n866 1
C_866   n867 0      1f

R_867   n868 n867 1
C_867   n868 0      1f

R_868   n869 n868 1
C_868   n869 0      1f

R_869   n870 n869 1
C_869   n870 0      1f

R_870   n871 n870 1
C_870   n871 0      1f

R_871   n872 n871 1
C_871   n872 0      1f

R_872   n873 n872 1
C_872   n873 0      1f

R_873   n874 n873 1
C_873   n874 0      1f

R_874   n875 n874 1
C_874   n875 0      1f

R_875   n876 n875 1
C_875   n876 0      1f

R_876   n877 n876 1
C_876   n877 0      1f

R_877   n878 n877 1
C_877   n878 0      1f

R_878   n879 n878 1
C_878   n879 0      1f

R_879   n880 n879 1
C_879   n880 0      1f

R_880   n881 n880 1
C_880   n881 0      1f

R_881   n882 n881 1
C_881   n882 0      1f

R_882   n883 n882 1
C_882   n883 0      1f

R_883   n884 n883 1
C_883   n884 0      1f

R_884   n885 n884 1
C_884   n885 0      1f

R_885   n886 n885 1
C_885   n886 0      1f

R_886   n887 n886 1
C_886   n887 0      1f

R_887   n888 n887 1
C_887   n888 0      1f

R_888   n889 n888 1
C_888   n889 0      1f

R_889   n890 n889 1
C_889   n890 0      1f

R_890   n891 n890 1
C_890   n891 0      1f

R_891   n892 n891 1
C_891   n892 0      1f

R_892   n893 n892 1
C_892   n893 0      1f

R_893   n894 n893 1
C_893   n894 0      1f

R_894   n895 n894 1
C_894   n895 0      1f

R_895   n896 n895 1
C_895   n896 0      1f

R_896   n897 n896 1
C_896   n897 0      1f

R_897   n898 n897 1
C_897   n898 0      1f

R_898   n899 n898 1
C_898   n899 0      1f

R_899   n900 n899 1
C_899   n900 0      1f

R_900   n901 n900 1
C_900   n901 0      1f

R_901   n902 n901 1
C_901   n902 0      1f

R_902   n903 n902 1
C_902   n903 0      1f

R_903   n904 n903 1
C_903   n904 0      1f

R_904   n905 n904 1
C_904   n905 0      1f

R_905   n906 n905 1
C_905   n906 0      1f

R_906   n907 n906 1
C_906   n907 0      1f

R_907   n908 n907 1
C_907   n908 0      1f

R_908   n909 n908 1
C_908   n909 0      1f

R_909   n910 n909 1
C_909   n910 0      1f

R_910   n911 n910 1
C_910   n911 0      1f

R_911   n912 n911 1
C_911   n912 0      1f

R_912   n913 n912 1
C_912   n913 0      1f

R_913   n914 n913 1
C_913   n914 0      1f

R_914   n915 n914 1
C_914   n915 0      1f

R_915   n916 n915 1
C_915   n916 0      1f

R_916   n917 n916 1
C_916   n917 0      1f

R_917   n918 n917 1
C_917   n918 0      1f

R_918   n919 n918 1
C_918   n919 0      1f

R_919   n920 n919 1
C_919   n920 0      1f

R_920   n921 n920 1
C_920   n921 0      1f

R_921   n922 n921 1
C_921   n922 0      1f

R_922   n923 n922 1
C_922   n923 0      1f

R_923   n924 n923 1
C_923   n924 0      1f

R_924   n925 n924 1
C_924   n925 0      1f

R_925   n926 n925 1
C_925   n926 0      1f

R_926   n927 n926 1
C_926   n927 0      1f

R_927   n928 n927 1
C_927   n928 0      1f

R_928   n929 n928 1
C_928   n929 0      1f

R_929   n930 n929 1
C_929   n930 0      1f

R_930   n931 n930 1
C_930   n931 0      1f

R_931   n932 n931 1
C_931   n932 0      1f

R_932   n933 n932 1
C_932   n933 0      1f

R_933   n934 n933 1
C_933   n934 0      1f

R_934   n935 n934 1
C_934   n935 0      1f

R_935   n936 n935 1
C_935   n936 0      1f

R_936   n937 n936 1
C_936   n937 0      1f

R_937   n938 n937 1
C_937   n938 0      1f

R_938   n939 n938 1
C_938   n939 0      1f

R_939   n940 n939 1
C_939   n940 0      1f

R_940   n941 n940 1
C_940   n941 0      1f

R_941   n942 n941 1
C_941   n942 0      1f

R_942   n943 n942 1
C_942   n943 0      1f

R_943   n944 n943 1
C_943   n944 0      1f

R_944   n945 n944 1
C_944   n945 0      1f

R_945   n946 n945 1
C_945   n946 0      1f

R_946   n947 n946 1
C_946   n947 0      1f

R_947   n948 n947 1
C_947   n948 0      1f

R_948   n949 n948 1
C_948   n949 0      1f

R_949   n950 n949 1
C_949   n950 0      1f

R_950   n951 n950 1
C_950   n951 0      1f

R_951   n952 n951 1
C_951   n952 0      1f

R_952   n953 n952 1
C_952   n953 0      1f

R_953   n954 n953 1
C_953   n954 0      1f

R_954   n955 n954 1
C_954   n955 0      1f

R_955   n956 n955 1
C_955   n956 0      1f

R_956   n957 n956 1
C_956   n957 0      1f

R_957   n958 n957 1
C_957   n958 0      1f

R_958   n959 n958 1
C_958   n959 0      1f

R_959   n960 n959 1
C_959   n960 0      1f

R_960   n961 n960 1
C_960   n961 0      1f

R_961   n962 n961 1
C_961   n962 0      1f

R_962   n963 n962 1
C_962   n963 0      1f

R_963   n964 n963 1
C_963   n964 0      1f

R_964   n965 n964 1
C_964   n965 0      1f

R_965   n966 n965 1
C_965   n966 0      1f

R_966   n967 n966 1
C_966   n967 0      1f

R_967   n968 n967 1
C_967   n968 0      1f

R_968   n969 n968 1
C_968   n969 0      1f

R_969   n970 n969 1
C_969   n970 0      1f

R_970   n971 n970 1
C_970   n971 0      1f

R_971   n972 n971 1
C_971   n972 0      1f

R_972   n973 n972 1
C_972   n973 0      1f

R_973   n974 n973 1
C_973   n974 0      1f

R_974   n975 n974 1
C_974   n975 0      1f

R_975   n976 n975 1
C_975   n976 0      1f

R_976   n977 n976 1
C_976   n977 0      1f

R_977   n978 n977 1
C_977   n978 0      1f

R_978   n979 n978 1
C_978   n979 0      1f

R_979   n980 n979 1
C_979   n980 0      1f

R_980   n981 n980 1
C_980   n981 0      1f

R_981   n982 n981 1
C_981   n982 0      1f

R_982   n983 n982 1
C_982   n983 0      1f

R_983   n984 n983 1
C_983   n984 0      1f

R_984   n985 n984 1
C_984   n985 0      1f

R_985   n986 n985 1
C_985   n986 0      1f

R_986   n987 n986 1
C_986   n987 0      1f

R_987   n988 n987 1
C_987   n988 0      1f

R_988   n989 n988 1
C_988   n989 0      1f

R_989   n990 n989 1
C_989   n990 0      1f

R_990   n991 n990 1
C_990   n991 0      1f

R_991   n992 n991 1
C_991   n992 0      1f

R_992   n993 n992 1
C_992   n993 0      1f

R_993   n994 n993 1
C_993   n994 0      1f

R_994   n995 n994 1
C_994   n995 0      1f

R_995   n996 n995 1
C_995   n996 0      1f

R_996   n997 n996 1
C_996   n997 0      1f

R_997   n998 n997 1
C_997   n998 0      1f

R_998   n999 n998 1
C_998   n999 0      1f

R_999   n1000 n999 1
C_999   n1000 0      1f

R_1000   n1001 n1000 1
C_1000   n1001 0      1f


.end