
*****************
* Include files *
*****************
.include '../memristor_ieee.cir'

***********
* Options *
***********
.option method=gear
.option reltol=1e-5 abstol=1e-9


***********
* Circuit *
***********
Xmemristor_ieee npos nneg memristor_ieee

***********
* Sources *
***********
Vin npos nneg AC 1  SIN(0V 2V  10MHz)

***************
* Simulations *
***************
* Operating point
.op

* AC analysis
*.ac dec 100 1e0 1e11

* Transient analysis
.tran 1e-9 1e-4

**********
* Output *
**********
.probe I V

.end

